//////////////////////////////////////////////////////////////////////////////////
// Module Name: image_gen
// Description: Generates a 46x46 pixel sprite/icon at coordinates (400, 400)
//////////////////////////////////////////////////////////////////////////////////

module image_gen #(
    parameter PIXELS_Y = 600,
    parameter PIXELS_X = 800
)(
    input  wire        clk,
    input  wire [31:0] row,   // Received as 32-bit vector from topmod
    input  wire [31:0] col,   // Received as 32-bit vector from topmod
	 input  wire [23:0]  obj_color,
	 input  wire [23:0]  bkg_color,
    output reg  [7:0]  red   = 8'h00,
    output reg  [7:0]  green = 8'h00,
    output reg  [7:0]  blue  = 8'h00
);

    // Sprite Data: 46 rows of 46-bit wide data
    reg [45:0] imageData [0:45];
    reg pixel_on;

    // Initialize the sprite data (replaces the VHDL constant array)
    initial begin
        imageData[0]  = 46'b0000000000000000001111111111000000000000000000;
        imageData[1]  = 46'b0000000000000111111111111111111110000000000000;
        imageData[2]  = 46'b0000000000001111111111111111111111000000000000;
        imageData[3]  = 46'b0000000000011111111111111111111111100000000000;
        imageData[4]  = 46'b0000000001111111111111111111111111111000000000;
        imageData[5]  = 46'b0000000011111111111111111111111111111100000000;
        imageData[6]  = 46'b0000001111111111111111111111111111111111000000;
        imageData[7]  = 46'b0000011111111111111111111111111111111111100000;
        imageData[8]  = 46'b0000111111111111111111111111111111111111110000;
        imageData[9]  = 46'b0000111111111111111111111111111111111111110000;
        imageData[10] = 46'b0001111111111111111111111111111111111111111000;
        imageData[11] = 46'b0001111111111111111111111111111111111111111000;
        imageData[12] = 46'b0011111111111111111111111111111111111111111100;
        imageData[13] = 46'b0111111111111100001111111111000011111111111110;
        imageData[14] = 46'b0111111111111000000111111110000001111111111110;
        imageData[15] = 46'b0111111111111000000111111110000001111111111110;
        imageData[16] = 46'b0111111111111000000111111110000001111111111110;
        imageData[17] = 46'b0111111111111000000111111110000001111111111110;
        imageData[18] = 46'b1111111111111100001111111111000011111111111111;
        imageData[19] = 46'b1111111111111111111111111111111111111111111111;
        imageData[20] = 46'b1111111111111111111111111111111111111111111111;
        imageData[21] = 46'b1111111111111111111111111111111111111111111111;
        imageData[22] = 46'b1111111111111111111111111111111111111111111111;
        imageData[23] = 46'b1111111111111111111111111111111111111111111111;
        imageData[24] = 46'b1111111111111111111111111111111111111111111111;
        imageData[25] = 46'b1111111111111111111111111111111111111111111111;
        imageData[26] = 46'b1111111111111111111111111111111111111111111111;
        imageData[27] = 46'b1111111111110000000000000000000000111111111111;
        imageData[28] = 46'b0111111111110000000000000000000000111111111110;
        imageData[29] = 46'b0111111111110000000000000000000000111111111110;
        imageData[30] = 46'b0111111111110000000000000000000000111111111110;
        imageData[31] = 46'b0111111111111000000000000000000001111111111110;
        imageData[32] = 46'b0111111111111000000000000000000001111111111110;
        imageData[33] = 46'b0011111111111100000000000000000011111111111100;
        imageData[34] = 46'b0001111111111100000000000000000011111111111000;
        imageData[35] = 46'b0001111111111111000000000000001111111111111000;
        imageData[36] = 46'b0000111111111111110000000000111111111111110000;
        imageData[37] = 46'b0000011111111111111000000001111111111111100000;
        imageData[38] = 46'b0000011111111111111111111111111111111111100000;
        imageData[39] = 46'b0000000111111111111111111111111111111110000000;
        imageData[40] = 46'b0000000011111111111111111111111111111100000000;
        imageData[41] = 46'b0000000001111111111111111111111111111000000000;
        imageData[42] = 46'b0000000000011111111111111111111111100000000000;
        imageData[43] = 46'b0000000000001111111111111111111111000000000000;
        imageData[44] = 46'b0000000000000011111111111111111100000000000000;
        imageData[45] = 46'b0000000000000000001111111111000000000000000000;
    end

   // Generation Logic
	always @(posedge clk) begin
		 if ((col >= 400 && col <= 445) && (row >= 400 && row <= 445)) begin
			  
			  pixel_on <= imageData[row-400][45-(col-400)];

			  if (pixel_on) begin
					red   <= obj_color[23:16];
					green <= obj_color[15:8];
					blue  <= obj_color[7:0];
			  end else begin
					// Pixel is inside the box, but part of the sprite background
					red   <= bkg_color[23:16];
					green <= bkg_color[15:8];
					blue  <= bkg_color[7:0];
			  end
			  
		 end else begin
			  // Entirely outside the 46x46 sprite box
			  red   <= 8'h00;
			  green <= 8'h00;
			  blue  <= 8'h00;
		 end
	end

endmodule